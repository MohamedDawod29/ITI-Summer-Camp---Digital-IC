Risc V architecture

Control Unit 
Extend Block     done
PCTarget       done